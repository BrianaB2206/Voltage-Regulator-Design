** Profile: "SCHEMATIC1-AC"  [ c:\users\brian\desktop\proiect1_simulation_files_boeru\schematics\proiect1_boeru-pspicefiles\schematic1\ac.sim ] 

** Creating circuit file "AC.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Users/brian/Desktop/V_regulator_Andreea/New folder/Lib_ModelePSpice_Anexa_1_a (1)/Modele_A1_lib/BC856B.lib" 
.LIB "C:/Users/brian/Desktop/V_regulator_Andreea/New folder/Lib_ModelePSpice_Anexa_1_a (1)/Modele_A1_lib/BC846B.lib" 
.LIB "C:/Users/brian/Desktop/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/THT/BC546.lib" 
.LIB "C:/Users/brian/Desktop/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/THT/TIP32C.LIB" 
.LIB "C:/Users/brian/Desktop/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/BZX84C2V7.lib" 
.LIB "C:/Users/brian/Desktop/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/MJD32CG.lib" 
.LIB "C:/Users/brian/Desktop/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/BC856B.lib" 
.LIB "C:/Users/brian/Desktop/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/BC846B.lib" 
.LIB "C:/Users/brian/Desktop/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/BZX84C5V1.lib" 
.LIB "C:/Users/brian/Desktop/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/BZX84C6V8.lib" 
* From [PSPICE NETLIST] section of C:\Users\brian\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
