** Profile: "SCHEMATIC1-Proiect1_Boeru_Bias"  [ E:\Proiect1_Boeru-PSpiceFiles\SCHEMATIC1\Proiect1_Boeru_Bias.sim ] 

** Creating circuit file "Proiect1_Boeru_Bias.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Users/brian/Desktop/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/MJD32CG.lib" 
.LIB "C:/Users/brian/Desktop/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/BC856B.lib" 
.LIB "C:/Users/brian/Desktop/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/BC846B.lib" 
.LIB "C:/Users/brian/Desktop/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/BZX84C5V1.lib" 
.LIB "C:/Users/brian/Desktop/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/BZX84C6V8.lib" 
* From [PSPICE NETLIST] section of C:\Users\brian\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
